module or_struct(a,b,o);

input a,b;
output o;

or(o,a,b);
endmodule