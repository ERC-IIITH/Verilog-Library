module xor_struct(a, b, o);

input a, b;
output o;

xor(o, a, b);

endmodule