module nand_struct(a, b, o);

input a, b;
output o;

nand(o, a, b);

endmodule