`timescale 1ns/1ps

module half_adder_struct
( output cout,sum,
  input a,b
  );
  
  
and a1(cout,a,b);
xor x1(sum,a,b);


endmodule
