module and_struct(a,b,o);

input a,b;
output o;

and(o,a,b);
endmodule